module out_mux();
